library IEEE;
use IEEE.std_logic_1164.all;

-- Package Declaration Section
package array_2D32bit is
 
  type Array2D is array (31 downto 0) of std_logic_vector(31 downto 0);

 
end package array_2D32bit;